library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity spi_master is
   generic (
      WTIME    : integer   := 100;
      TXBITS   : integer   := 16;
      RXBITS   : integer   := 8
      );
   port ( 
      clock    : in  std_logic;
      reset    : in  std_logic;
      txd      : in  std_logic_vector(TXBITS-1 downto 0);
      rxd      : out std_logic_vector(RXBITS-1 downto 0);
      start    : in  std_logic;
      ready    : out std_logic;
      miso     : in  std_logic;
      mosi     : out std_logic;
      sclk     : out std_logic;
      cs       : out std_logic
      );
end spi_master;

architecture Behavioral of spi_master is

----------------------------------------
------  WRITE YOUR CODE HERE  ----------
----------------------------------------
   
begin

----------------------------------------
------  WRITE YOUR CODE HERE  ----------
-- and delete the following 3 lines  ---
----------------------------------------   
cs <= '1'; 
sclk <= '0';
mosi <= miso; 

end Behavioral;

